magic
tech sky130A
magscale 1 2
timestamp 1729232797
<< psubdiff >>
rect 1081 585 1180 619
rect 2280 585 2363 619
rect 1081 504 1115 585
rect 2329 504 2363 585
rect 1081 -163 1115 -130
rect 2329 -163 2363 -130
rect 1081 -197 1180 -163
rect 2280 -197 2363 -163
<< psubdiffcont >>
rect 1180 585 2280 619
rect 1081 -130 1115 504
rect 2329 -130 2363 504
rect 1180 -197 2280 -163
<< poly >>
rect 1165 538 1257 554
rect 1165 504 1181 538
rect 1215 504 1257 538
rect 1165 488 1257 504
rect 1227 466 1257 488
rect 2187 538 2279 554
rect 2187 504 2229 538
rect 2263 504 2279 538
rect 2187 488 2279 504
rect 2187 462 2217 488
rect 1227 -66 1257 -44
rect 1165 -82 1257 -66
rect 1165 -116 1181 -82
rect 1215 -116 1257 -82
rect 1165 -132 1257 -116
rect 2187 -66 2217 -15
rect 2187 -82 2279 -66
rect 2187 -116 2229 -82
rect 2263 -116 2279 -82
rect 2187 -132 2279 -116
<< polycont >>
rect 1181 504 1215 538
rect 2229 504 2263 538
rect 1181 -116 1215 -82
rect 2229 -116 2263 -82
<< locali >>
rect 1081 585 1180 619
rect 2280 585 2363 619
rect 1081 504 1115 585
rect 1165 504 1181 538
rect 1215 504 1231 538
rect 2213 504 2229 538
rect 2263 504 2279 538
rect 2329 504 2363 585
rect 1181 466 1215 504
rect 2229 462 2263 504
rect 1181 -82 1215 -44
rect 2229 -82 2263 -15
rect 1165 -116 1181 -82
rect 1215 -116 1231 -82
rect 2213 -116 2229 -82
rect 2263 -116 2279 -82
rect 1081 -163 1115 -130
rect 2329 -163 2363 -130
rect 1081 -197 1180 -163
rect 2280 -197 2363 -163
<< viali >>
rect 1487 585 1521 619
rect 1923 585 1957 619
rect 1181 504 1215 538
rect 2229 504 2263 538
rect 1181 -116 1215 -82
rect 2229 -116 2263 -82
rect 1487 -197 1521 -163
rect 1923 -197 1957 -163
<< metal1 >>
rect 1468 576 1478 628
rect 1530 576 1540 628
rect 1904 576 1914 628
rect 1966 576 1976 628
rect 1169 538 1227 544
rect 1169 504 1181 538
rect 1215 504 1227 538
rect 1169 498 1227 504
rect 2217 538 2275 544
rect 2217 504 2229 538
rect 2263 504 2275 538
rect 2217 498 2275 504
rect 1175 466 1221 498
rect 2223 466 2269 498
rect 1175 266 1309 466
rect 1468 277 1478 453
rect 1530 277 1540 453
rect 1686 278 1696 454
rect 1748 278 1758 454
rect 1904 278 1914 454
rect 1966 278 1976 454
rect 2135 266 2269 466
rect 1262 234 1308 266
rect 2135 234 2181 266
rect 1262 188 2181 234
rect 1262 187 2125 188
rect 1175 144 1309 156
rect 1175 -31 1260 144
rect 1175 -44 1213 -31
rect 1219 -32 1260 -31
rect 1312 -32 1322 144
rect 1468 -32 1478 144
rect 1530 -32 1540 144
rect 1219 -44 1309 -32
rect 1699 -44 1745 187
rect 2135 144 2269 156
rect 1904 -32 1914 144
rect 1966 -32 1976 144
rect 2122 -32 2132 144
rect 2184 -32 2269 144
rect 2135 -44 2269 -32
rect 1175 -76 1221 -44
rect 2223 -76 2269 -44
rect 1169 -82 1227 -76
rect 1169 -116 1181 -82
rect 1215 -116 1227 -82
rect 1169 -122 1227 -116
rect 2217 -82 2275 -76
rect 2217 -116 2229 -82
rect 2263 -116 2275 -82
rect 2217 -122 2275 -116
rect 1468 -206 1478 -154
rect 1530 -206 1540 -154
rect 1904 -206 1914 -154
rect 1966 -206 1976 -154
<< via1 >>
rect 1478 619 1530 628
rect 1478 585 1487 619
rect 1487 585 1521 619
rect 1521 585 1530 619
rect 1478 576 1530 585
rect 1914 619 1966 628
rect 1914 585 1923 619
rect 1923 585 1957 619
rect 1957 585 1966 619
rect 1914 576 1966 585
rect 1478 277 1530 453
rect 1696 278 1748 454
rect 1914 278 1966 454
rect 1260 -32 1312 144
rect 1478 -32 1530 144
rect 1914 -32 1966 144
rect 2132 -32 2184 144
rect 1478 -163 1530 -154
rect 1478 -197 1487 -163
rect 1487 -197 1521 -163
rect 1521 -197 1530 -163
rect 1478 -206 1530 -197
rect 1914 -163 1966 -154
rect 1914 -197 1923 -163
rect 1923 -197 1957 -163
rect 1957 -197 1966 -163
rect 1914 -206 1966 -197
<< metal2 >>
rect 1478 628 1530 638
rect 1478 453 1530 576
rect 1914 628 1966 638
rect 1478 267 1530 277
rect 1696 454 1748 464
rect 1696 237 1748 278
rect 1914 454 1966 576
rect 1914 268 1966 278
rect 1260 185 2184 237
rect 1260 144 1312 185
rect 1260 -42 1312 -32
rect 1478 144 1530 154
rect 1478 -154 1530 -32
rect 1478 -216 1530 -206
rect 1914 144 1966 154
rect 1914 -154 1966 -32
rect 2132 144 2184 185
rect 2132 -42 2184 -32
rect 1914 -216 1966 -206
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729220960
transform 1 0 2202 0 1 56
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729220960
transform 1 0 1242 0 1 56
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729220960
transform 1 0 1242 0 1 366
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729220960
transform 1 0 2202 0 1 366
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_YJHC9X  sky130_fd_pr__nfet_01v8_YJHC9X_0
timestamp 1729231875
transform 1 0 1722 0 1 211
box -465 -343 465 343
<< labels >>
flabel metal1 1248 383 1248 383 0 FreeSans 480 0 0 0 d8
port 1 nsew
flabel metal1 1243 49 1243 49 0 FreeSans 480 0 0 0 d9
port 2 nsew
flabel locali 2292 609 2292 609 0 FreeSans 480 0 0 0 gnd
port 0 nsew
<< end >>
