magic
tech sky130A
magscale 1 2
timestamp 1729433138
<< locali >>
rect 1046 3790 1134 3824
<< viali >>
rect 1012 3790 1046 3824
<< metal1 >>
rect -30 4161 140 4195
rect -30 1568 6 4161
rect 1000 3824 1135 3833
rect 1000 3790 1012 3824
rect 1046 3790 1135 3824
rect 1000 3781 1135 3790
rect 1255 3039 1265 3091
rect 1441 3039 1451 3091
rect 1565 3036 1575 3088
rect 1751 3036 1761 3088
rect 786 2836 1156 2882
rect 304 2753 314 2805
rect 366 2753 376 2805
rect 1417 1768 1451 1891
rect -30 1534 140 1568
<< via1 >>
rect 1265 3039 1441 3091
rect 1575 3036 1751 3088
rect 314 2753 366 2805
<< metal2 >>
rect 1265 3091 1441 3101
rect 314 2805 366 3076
rect 1265 2829 1441 3039
rect 1265 2763 1441 2773
rect 1575 3088 1751 3098
rect 1575 3026 1751 3036
rect 314 2743 366 2753
rect 1575 2268 1627 3026
rect 1242 1817 1310 1891
rect 786 442 844 444
rect 1327 442 1383 452
rect 786 386 1327 442
rect 1383 386 1392 442
rect 786 367 844 386
rect 1327 376 1383 386
<< via2 >>
rect 1265 2773 1441 2829
rect 1327 386 1383 442
<< metal3 >>
rect 547 3584 619 3735
rect 1255 2829 1451 2834
rect 1255 2773 1265 2829
rect 1441 2773 1451 2829
rect 1255 2768 1451 2773
rect 1317 442 1393 712
rect 1317 386 1327 442
rect 1383 386 1393 442
rect 1317 381 1393 386
use nmoscs2  nmoscs2_0
timestamp 1729232797
transform 0 -1 1719 1 0 1867
box 1081 -216 2363 638
use nmoscs  nmoscs_0
timestamp 1729186456
transform 1 0 183 0 1 4165
box -213 -1253 899 151
use pmoscs  pmoscs_0
timestamp 1729152905
transform 1 0 148 0 1 752
box -178 -740 820 2160
use pmosdiff  pmosdiff_0
timestamp 1729428050
transform 1 0 1054 0 1 684
box -98 -671 700 2228
<< labels >>
flabel viali 1025 3807 1025 3807 0 FreeSans 480 0 0 0 gnd
port 1 nsew
flabel metal1 818 2856 818 2856 0 FreeSans 480 0 0 0 vdd
port 0 nsew
flabel metal2 1592 2680 1592 2680 0 FreeSans 480 0 0 0 out
port 2 nsew
flabel metal2 1275 1841 1275 1841 0 FreeSans 480 0 0 0 vip
port 3 nsew
flabel metal1 1431 1833 1431 1833 0 FreeSans 480 0 0 0 vin
port 4 nsew
flabel metal3 583 3660 583 3660 0 FreeSans 480 0 0 0 rs
port 5 nsew
<< end >>
