magic
tech sky130A
magscale 1 2
timestamp 1729242668
<< error_p >>
rect -223 338 223 556
rect -223 18 223 236
rect -223 -302 223 -84
<< nwell >>
rect -223 338 223 622
rect -223 18 223 302
rect -223 -302 223 -18
rect -223 -622 223 -338
<< pmos >>
rect -129 438 -29 522
rect 29 438 129 522
rect -129 118 -29 202
rect 29 118 129 202
rect -129 -202 -29 -118
rect 29 -202 129 -118
rect -129 -522 -29 -438
rect 29 -522 129 -438
<< pdiff >>
rect -187 510 -129 522
rect -187 450 -175 510
rect -141 450 -129 510
rect -187 438 -129 450
rect -29 510 29 522
rect -29 450 -17 510
rect 17 450 29 510
rect -29 438 29 450
rect 129 510 187 522
rect 129 450 141 510
rect 175 450 187 510
rect 129 438 187 450
rect -187 190 -129 202
rect -187 130 -175 190
rect -141 130 -129 190
rect -187 118 -129 130
rect -29 190 29 202
rect -29 130 -17 190
rect 17 130 29 190
rect -29 118 29 130
rect 129 190 187 202
rect 129 130 141 190
rect 175 130 187 190
rect 129 118 187 130
rect -187 -130 -129 -118
rect -187 -190 -175 -130
rect -141 -190 -129 -130
rect -187 -202 -129 -190
rect -29 -130 29 -118
rect -29 -190 -17 -130
rect 17 -190 29 -130
rect -29 -202 29 -190
rect 129 -130 187 -118
rect 129 -190 141 -130
rect 175 -190 187 -130
rect 129 -202 187 -190
rect -187 -450 -129 -438
rect -187 -510 -175 -450
rect -141 -510 -129 -450
rect -187 -522 -129 -510
rect -29 -450 29 -438
rect -29 -510 -17 -450
rect 17 -510 29 -450
rect -29 -522 29 -510
rect 129 -450 187 -438
rect 129 -510 141 -450
rect 175 -510 187 -450
rect 129 -522 187 -510
<< pdiffc >>
rect -175 450 -141 510
rect -17 450 17 510
rect 141 450 175 510
rect -175 130 -141 190
rect -17 130 17 190
rect 141 130 175 190
rect -175 -190 -141 -130
rect -17 -190 17 -130
rect 141 -190 175 -130
rect -175 -510 -141 -450
rect -17 -510 17 -450
rect 141 -510 175 -450
<< poly >>
rect -129 603 -29 619
rect -129 569 -113 603
rect -45 569 -29 603
rect -129 522 -29 569
rect 29 603 129 619
rect 29 569 45 603
rect 113 569 129 603
rect 29 522 129 569
rect -129 391 -29 438
rect -129 357 -113 391
rect -45 357 -29 391
rect -129 341 -29 357
rect 29 391 129 438
rect 29 357 45 391
rect 113 357 129 391
rect 29 341 129 357
rect -129 283 -29 299
rect -129 249 -113 283
rect -45 249 -29 283
rect -129 202 -29 249
rect 29 283 129 299
rect 29 249 45 283
rect 113 249 129 283
rect 29 202 129 249
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect -129 -249 -29 -202
rect -129 -283 -113 -249
rect -45 -283 -29 -249
rect -129 -299 -29 -283
rect 29 -249 129 -202
rect 29 -283 45 -249
rect 113 -283 129 -249
rect 29 -299 129 -283
rect -129 -357 -29 -341
rect -129 -391 -113 -357
rect -45 -391 -29 -357
rect -129 -438 -29 -391
rect 29 -357 129 -341
rect 29 -391 45 -357
rect 113 -391 129 -357
rect 29 -438 129 -391
rect -129 -569 -29 -522
rect -129 -603 -113 -569
rect -45 -603 -29 -569
rect -129 -619 -29 -603
rect 29 -569 129 -522
rect 29 -603 45 -569
rect 113 -603 129 -569
rect 29 -619 129 -603
<< polycont >>
rect -113 569 -45 603
rect 45 569 113 603
rect -113 357 -45 391
rect 45 357 113 391
rect -113 249 -45 283
rect 45 249 113 283
rect -113 37 -45 71
rect 45 37 113 71
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -113 -283 -45 -249
rect 45 -283 113 -249
rect -113 -391 -45 -357
rect 45 -391 113 -357
rect -113 -603 -45 -569
rect 45 -603 113 -569
<< locali >>
rect -129 569 -113 603
rect -45 569 -29 603
rect 29 569 45 603
rect 113 569 129 603
rect -175 510 -141 526
rect -175 434 -141 450
rect -17 510 17 526
rect -17 434 17 450
rect 141 510 175 526
rect 141 434 175 450
rect -129 357 -113 391
rect -45 357 -29 391
rect 29 357 45 391
rect 113 357 129 391
rect -129 249 -113 283
rect -45 249 -29 283
rect 29 249 45 283
rect 113 249 129 283
rect -175 190 -141 206
rect -175 114 -141 130
rect -17 190 17 206
rect -17 114 17 130
rect 141 190 175 206
rect 141 114 175 130
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect -175 -130 -141 -114
rect -175 -206 -141 -190
rect -17 -130 17 -114
rect -17 -206 17 -190
rect 141 -130 175 -114
rect 141 -206 175 -190
rect -129 -283 -113 -249
rect -45 -283 -29 -249
rect 29 -283 45 -249
rect 113 -283 129 -249
rect -129 -391 -113 -357
rect -45 -391 -29 -357
rect 29 -391 45 -357
rect 113 -391 129 -357
rect -175 -450 -141 -434
rect -175 -526 -141 -510
rect -17 -450 17 -434
rect -17 -526 17 -510
rect 141 -450 175 -434
rect 141 -526 175 -510
rect -129 -603 -113 -569
rect -45 -603 -29 -569
rect 29 -603 45 -569
rect 113 -603 129 -569
<< viali >>
rect -113 569 -45 603
rect 45 569 113 603
rect -175 450 -141 510
rect -17 450 17 510
rect 141 450 175 510
rect -113 357 -45 391
rect 45 357 113 391
rect -113 249 -45 283
rect 45 249 113 283
rect -175 130 -141 190
rect -17 130 17 190
rect 141 130 175 190
rect -113 37 -45 71
rect 45 37 113 71
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect -175 -190 -141 -130
rect -17 -190 17 -130
rect 141 -190 175 -130
rect -113 -283 -45 -249
rect 45 -283 113 -249
rect -113 -391 -45 -357
rect 45 -391 113 -357
rect -175 -510 -141 -450
rect -17 -510 17 -450
rect 141 -510 175 -450
rect -113 -603 -45 -569
rect 45 -603 113 -569
<< metal1 >>
rect -125 603 -33 609
rect -125 569 -113 603
rect -45 569 -33 603
rect -125 563 -33 569
rect 33 603 125 609
rect 33 569 45 603
rect 113 569 125 603
rect 33 563 125 569
rect -181 510 -135 522
rect -181 450 -175 510
rect -141 450 -135 510
rect -181 438 -135 450
rect -23 510 23 522
rect -23 450 -17 510
rect 17 450 23 510
rect -23 438 23 450
rect 135 510 181 522
rect 135 450 141 510
rect 175 450 181 510
rect 135 438 181 450
rect -125 391 -33 397
rect -125 357 -113 391
rect -45 357 -33 391
rect -125 351 -33 357
rect 33 391 125 397
rect 33 357 45 391
rect 113 357 125 391
rect 33 351 125 357
rect -125 283 -33 289
rect -125 249 -113 283
rect -45 249 -33 283
rect -125 243 -33 249
rect 33 283 125 289
rect 33 249 45 283
rect 113 249 125 283
rect 33 243 125 249
rect -181 190 -135 202
rect -181 130 -175 190
rect -141 130 -135 190
rect -181 118 -135 130
rect -23 190 23 202
rect -23 130 -17 190
rect 17 130 23 190
rect -23 118 23 130
rect 135 190 181 202
rect 135 130 141 190
rect 175 130 181 190
rect 135 118 181 130
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect -181 -130 -135 -118
rect -181 -190 -175 -130
rect -141 -190 -135 -130
rect -181 -202 -135 -190
rect -23 -130 23 -118
rect -23 -190 -17 -130
rect 17 -190 23 -130
rect -23 -202 23 -190
rect 135 -130 181 -118
rect 135 -190 141 -130
rect 175 -190 181 -130
rect 135 -202 181 -190
rect -125 -249 -33 -243
rect -125 -283 -113 -249
rect -45 -283 -33 -249
rect -125 -289 -33 -283
rect 33 -249 125 -243
rect 33 -283 45 -249
rect 113 -283 125 -249
rect 33 -289 125 -283
rect -125 -357 -33 -351
rect -125 -391 -113 -357
rect -45 -391 -33 -357
rect -125 -397 -33 -391
rect 33 -357 125 -351
rect 33 -391 45 -357
rect 113 -391 125 -357
rect 33 -397 125 -391
rect -181 -450 -135 -438
rect -181 -510 -175 -450
rect -141 -510 -135 -450
rect -181 -522 -135 -510
rect -23 -450 23 -438
rect -23 -510 -17 -450
rect 17 -510 23 -450
rect -23 -522 23 -510
rect 135 -450 181 -438
rect 135 -510 141 -450
rect 175 -510 181 -450
rect 135 -522 181 -510
rect -125 -569 -33 -563
rect -125 -603 -113 -569
rect -45 -603 -33 -569
rect -125 -609 -33 -603
rect 33 -569 125 -563
rect 33 -603 45 -569
rect 113 -603 125 -569
rect 33 -609 125 -603
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.5 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
