magic
tech sky130A
magscale 1 2
timestamp 1729186456
<< pwell >>
rect -213 -1253 899 151
<< psubdiff >>
rect -177 81 263 115
rect 421 81 863 115
rect -177 -427 -143 81
rect -177 -1183 -143 -667
rect 829 -427 863 81
rect 829 -1183 863 -667
rect -177 -1217 263 -1183
rect 421 -1217 863 -1183
<< psubdiffcont >>
rect 263 81 421 115
rect -177 -667 -143 -427
rect 829 -667 863 -427
rect 263 -1217 421 -1183
<< poly >>
rect -93 30 -1 46
rect -93 -4 -77 30
rect -43 -4 -1 30
rect -93 -20 -1 -4
rect -31 -42 -1 -20
rect 687 30 779 46
rect 687 -4 729 30
rect 763 -4 779 30
rect 687 -20 779 -4
rect 687 -42 717 -20
rect -31 -1082 -1 -1060
rect -93 -1098 -1 -1082
rect -93 -1132 -77 -1098
rect -43 -1132 -1 -1098
rect -93 -1148 -1 -1132
rect 687 -1082 717 -1080
rect 687 -1098 779 -1082
rect 687 -1132 729 -1098
rect 763 -1132 779 -1098
rect 687 -1148 779 -1132
<< polycont >>
rect -77 -4 -43 30
rect 729 -4 763 30
rect -77 -1132 -43 -1098
rect 729 -1132 763 -1098
<< locali >>
rect -177 81 263 115
rect 421 81 863 115
rect -177 -427 -143 81
rect -93 -4 -77 30
rect -43 -4 -27 30
rect -77 -42 -43 -4
rect 269 -39 303 81
rect 713 -4 729 30
rect 763 -4 779 30
rect 729 -42 763 -4
rect 829 -427 863 81
rect -177 -1183 -143 -667
rect -77 -1098 -43 -1060
rect -93 -1132 -77 -1098
rect -43 -1132 -27 -1098
rect 383 -1183 417 -1048
rect 729 -1098 763 -1060
rect 713 -1132 729 -1098
rect 763 -1132 779 -1098
rect 829 -1183 863 -667
rect -177 -1217 263 -1183
rect 421 -1217 863 -1183
<< viali >>
rect 269 81 303 115
rect -77 -4 -43 30
rect 729 -4 763 30
rect 269 -430 303 -54
rect 383 -430 417 -54
rect 269 -1048 303 -672
rect 383 -1048 417 -672
rect -77 -1132 -43 -1098
rect 729 -1132 763 -1098
rect 383 -1217 417 -1183
<< metal1 >>
rect 257 115 315 121
rect 257 81 269 115
rect 303 81 315 115
rect 257 75 315 81
rect -89 30 -31 36
rect -89 -4 -77 30
rect -43 -4 -31 30
rect -89 -10 -31 -4
rect -83 -42 -37 -10
rect -83 -442 51 -42
rect 263 -54 309 75
rect 717 30 775 36
rect 717 -4 729 30
rect 763 -4 775 30
rect 717 -10 775 -4
rect 723 -42 769 -10
rect 377 -54 423 -42
rect 635 -54 769 -42
rect 250 -430 260 -54
rect 312 -430 322 -54
rect 364 -430 374 -54
rect 426 -430 436 -54
rect 622 -430 632 -54
rect 684 -430 769 -54
rect 263 -442 309 -430
rect 377 -442 423 -430
rect 635 -442 769 -430
rect 5 -474 51 -442
rect 5 -530 625 -474
rect 5 -572 681 -530
rect 61 -628 681 -572
rect 635 -660 681 -628
rect -83 -672 51 -660
rect 263 -672 309 -660
rect 377 -672 423 -660
rect -83 -1048 2 -672
rect 54 -1048 64 -672
rect 250 -1048 260 -672
rect 312 -1048 322 -672
rect 364 -1048 374 -672
rect 426 -1048 436 -672
rect -83 -1060 51 -1048
rect 263 -1060 309 -1048
rect -83 -1092 -37 -1060
rect -89 -1098 -31 -1092
rect -89 -1132 -77 -1098
rect -43 -1132 -31 -1098
rect -89 -1138 -31 -1132
rect 374 -1177 426 -1048
rect 635 -1060 769 -660
rect 723 -1092 769 -1060
rect 717 -1098 775 -1092
rect 717 -1132 729 -1098
rect 763 -1132 775 -1098
rect 717 -1138 775 -1132
rect 371 -1183 429 -1177
rect 371 -1217 383 -1183
rect 417 -1217 429 -1183
rect 371 -1223 429 -1217
<< via1 >>
rect 260 -430 269 -54
rect 269 -430 303 -54
rect 303 -430 312 -54
rect 374 -430 383 -54
rect 383 -430 417 -54
rect 417 -430 426 -54
rect 632 -430 684 -54
rect 2 -1048 54 -672
rect 260 -1048 269 -672
rect 269 -1048 303 -672
rect 303 -1048 312 -672
rect 374 -1048 383 -672
rect 383 -1048 417 -672
rect 417 -1048 426 -672
<< metal2 >>
rect 1 -13 684 39
rect 2 -672 54 -13
rect 260 -54 312 -48
rect 260 -440 312 -430
rect 372 -54 428 -44
rect 372 -440 428 -430
rect 632 -54 684 -13
rect 263 -530 309 -440
rect 263 -572 423 -530
rect 377 -662 423 -572
rect 2 -1089 54 -1048
rect 258 -672 314 -662
rect 258 -1058 314 -1048
rect 374 -672 426 -662
rect 374 -1060 426 -1048
rect 632 -1089 684 -430
rect 2 -1141 684 -1089
<< via2 >>
rect 372 -430 374 -54
rect 374 -430 426 -54
rect 426 -430 428 -54
rect 258 -1048 260 -672
rect 260 -1048 312 -672
rect 312 -1048 314 -672
<< metal3 >>
rect 362 -54 438 -49
rect 358 -430 372 -54
rect 428 -430 442 -54
rect 362 -435 438 -430
rect 364 -521 436 -435
rect 250 -581 436 -521
rect 250 -667 322 -581
rect 248 -672 324 -667
rect 244 -1048 258 -672
rect 314 -1048 328 -672
rect 248 -1053 324 -1048
use sky130_fd_pr__nfet_01v8_27FZYL  sky130_fd_pr__nfet_01v8_27FZYL_0
timestamp 1729158022
transform 1 0 343 0 1 -273
box -344 -257 344 257
use sky130_fd_pr__nfet_01v8_Q6296P  sky130_fd_pr__nfet_01v8_Q6296P_0
timestamp 1729158022
transform 1 0 343 0 1 -829
box -344 -257 344 257
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_0
timestamp 1729171183
transform 1 0 702 0 1 -860
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_1
timestamp 1729171183
transform 1 0 -16 0 1 -242
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_2
timestamp 1729171183
transform 1 0 -16 0 1 -860
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_3
timestamp 1729171183
transform 1 0 702 0 1 -242
box -73 -226 73 226
<< labels >>
flabel viali 398 -1196 398 -1196 0 FreeSans 480 0 0 0 gnd
port 0 nsew
flabel metal1 -17 -169 -17 -169 0 FreeSans 480 0 0 0 d3
port 1 nsew
flabel metal2 653 -12 653 -12 0 FreeSans 480 0 0 0 d4
port 2 nsew
flabel metal3 395 -462 395 -462 0 FreeSans 480 0 0 0 rs
port 3 nsew
<< end >>
