magic
tech sky130A
magscale 1 2
timestamp 1729428050
<< nwell >>
rect -98 -671 700 2228
<< pmos >>
rect 488 220 518 221
<< pdiff >>
rect 518 220 576 221
<< nsubdiff >>
rect -62 2158 33 2192
rect 569 2158 664 2192
rect -62 1690 -28 2158
rect 630 1690 664 2158
rect -62 -600 -28 -132
rect 630 -600 664 -132
rect -62 -634 33 -600
rect 569 -634 664 -600
<< nsubdiffcont >>
rect 33 2158 569 2192
rect -62 -132 -28 1690
rect 630 -132 664 1690
rect 33 -634 569 -600
<< poly >>
rect 84 1306 114 1326
rect 22 1290 114 1306
rect 22 1256 38 1290
rect 72 1256 114 1290
rect 22 1240 114 1256
rect 488 1306 518 1322
rect 488 1290 580 1306
rect 488 1256 530 1290
rect 564 1256 580 1290
rect 488 1240 580 1256
rect 22 1124 114 1140
rect 22 1090 38 1124
rect 72 1090 114 1124
rect 22 1074 114 1090
rect 84 1051 114 1074
rect 488 1124 580 1140
rect 488 1090 530 1124
rect 564 1090 580 1124
rect 488 1074 580 1090
rect 488 1043 518 1074
rect 84 484 114 527
rect 22 468 114 484
rect 22 434 38 468
rect 72 434 114 468
rect 22 418 114 434
rect 488 484 518 500
rect 488 468 580 484
rect 488 434 530 468
rect 564 434 580 468
rect 488 418 580 434
rect 22 302 114 318
rect 22 268 38 302
rect 72 268 114 302
rect 22 252 114 268
rect 84 221 114 252
rect 488 302 580 318
rect 488 268 530 302
rect 564 268 580 302
rect 488 252 580 268
rect 488 221 518 252
<< polycont >>
rect 38 1256 72 1290
rect 530 1256 564 1290
rect 38 1090 72 1124
rect 530 1090 564 1124
rect 38 434 72 468
rect 530 434 564 468
rect 38 268 72 302
rect 530 268 564 302
<< locali >>
rect -62 2158 33 2192
rect 569 2158 664 2192
rect -62 1690 -28 2158
rect 630 1690 664 2158
rect 38 1290 72 1364
rect 530 1290 564 1354
rect 22 1256 38 1290
rect 72 1256 88 1290
rect 514 1256 530 1290
rect 564 1256 580 1290
rect 22 1090 38 1124
rect 72 1090 88 1124
rect 514 1090 530 1124
rect 564 1090 580 1124
rect 38 1043 72 1090
rect 530 1044 564 1090
rect 38 468 72 527
rect 530 468 564 512
rect 22 434 38 468
rect 72 434 88 468
rect 514 434 530 468
rect 564 434 580 468
rect 22 268 38 302
rect 72 268 88 302
rect 514 268 530 302
rect 564 268 580 302
rect 38 221 72 268
rect 530 220 564 268
rect -62 -600 -28 -132
rect 630 -600 664 -132
rect -62 -634 33 -600
rect 569 -634 664 -600
<< viali >>
rect 105 2158 497 2192
rect 38 1256 72 1290
rect 530 1256 564 1290
rect 38 1090 72 1124
rect 530 1090 564 1124
rect 38 434 72 468
rect 530 434 564 468
rect 38 268 72 302
rect 530 268 564 302
<< metal1 >>
rect 93 2192 509 2198
rect 93 2158 105 2192
rect 497 2158 509 2192
rect 93 2152 509 2158
rect 32 1525 166 1537
rect 436 1525 570 1537
rect 32 1349 117 1525
rect 169 1349 179 1525
rect 265 1349 275 1525
rect 327 1349 337 1525
rect 436 1349 521 1525
rect 573 1349 583 1525
rect 32 1337 166 1349
rect 436 1337 570 1349
rect 32 1296 78 1337
rect 26 1290 84 1296
rect 26 1256 38 1290
rect 72 1256 84 1290
rect 26 1250 84 1256
rect 205 1207 239 1290
rect 336 1247 346 1299
rect 414 1247 424 1299
rect 524 1296 570 1337
rect 518 1290 576 1296
rect 518 1256 530 1290
rect 564 1256 576 1290
rect 518 1250 576 1256
rect 205 1173 397 1207
rect 26 1124 84 1130
rect 26 1090 38 1124
rect 72 1090 84 1124
rect 26 1084 84 1090
rect 32 1043 77 1084
rect 178 1081 188 1133
rect 256 1081 266 1133
rect 363 1090 397 1173
rect 518 1124 576 1130
rect 518 1090 530 1124
rect 564 1090 576 1124
rect 518 1084 576 1090
rect 524 1043 570 1084
rect 32 1031 166 1043
rect 436 1031 570 1043
rect -16 855 29 1031
rect 81 855 166 1031
rect 265 855 275 1031
rect 327 855 337 1031
rect 423 855 433 1031
rect 485 855 570 1031
rect 32 843 166 855
rect 436 843 570 855
rect 32 703 166 715
rect 436 703 570 715
rect -16 527 29 703
rect 81 527 166 703
rect 265 527 275 703
rect 327 527 337 703
rect 423 527 433 703
rect 485 527 570 703
rect 32 515 166 527
rect 436 515 570 527
rect 32 474 77 515
rect 26 468 84 474
rect 26 434 38 468
rect 72 434 84 468
rect 26 428 84 434
rect 178 425 188 477
rect 256 425 266 477
rect 523 474 570 515
rect 518 468 576 474
rect 518 434 530 468
rect 564 434 576 468
rect 518 428 576 434
rect 363 385 397 428
rect 205 351 397 385
rect 205 308 239 351
rect 26 302 84 308
rect 26 268 38 302
rect 72 268 84 302
rect 26 262 84 268
rect 32 221 78 262
rect 336 259 346 311
rect 414 259 424 311
rect 518 302 576 308
rect 518 268 530 302
rect 564 268 576 302
rect 518 262 576 268
rect 524 221 570 262
rect 32 209 166 221
rect 436 209 570 221
rect 32 33 117 209
rect 169 33 179 209
rect 265 33 275 209
rect 327 33 337 209
rect 436 33 521 209
rect 573 33 583 209
rect 32 21 166 33
rect 436 21 570 33
<< via1 >>
rect 117 1349 169 1525
rect 275 1349 327 1525
rect 521 1349 573 1525
rect 346 1247 414 1299
rect 188 1081 256 1133
rect 29 855 81 1031
rect 275 855 327 1031
rect 433 855 485 1031
rect 29 527 81 703
rect 275 527 327 703
rect 433 527 485 703
rect 188 425 256 477
rect 346 259 414 311
rect 117 33 169 209
rect 275 33 327 209
rect 521 33 573 209
<< metal2 >>
rect 29 1585 573 1637
rect 29 1031 81 1585
rect 115 1525 171 1535
rect 115 1339 171 1349
rect 273 1525 329 1535
rect 273 1339 329 1349
rect 521 1525 573 1585
rect 275 1337 327 1339
rect 346 1299 414 1309
rect 346 1207 414 1247
rect 188 1173 414 1207
rect 188 1133 256 1173
rect 188 1071 256 1081
rect 275 1041 327 1043
rect 29 703 81 855
rect 273 1031 329 1041
rect 273 845 329 855
rect 431 1031 487 1041
rect 431 845 487 855
rect 275 713 327 845
rect 29 -27 81 527
rect 273 703 329 713
rect 273 517 329 527
rect 431 703 487 713
rect 431 517 487 527
rect 275 515 327 517
rect 188 477 256 487
rect 188 385 256 425
rect 188 351 414 385
rect 346 311 414 351
rect 346 249 414 259
rect 275 219 327 221
rect 115 209 171 219
rect 115 23 171 33
rect 273 209 329 219
rect 273 23 329 33
rect 521 209 573 1349
rect 521 -27 573 33
rect 29 -79 573 -27
<< via2 >>
rect 115 1349 117 1525
rect 117 1349 169 1525
rect 169 1349 171 1525
rect 273 1349 275 1525
rect 275 1349 327 1525
rect 327 1349 329 1525
rect 273 855 275 1031
rect 275 855 327 1031
rect 327 855 329 1031
rect 431 855 433 1031
rect 433 855 485 1031
rect 485 855 487 1031
rect 273 527 275 703
rect 275 527 327 703
rect 327 527 329 703
rect 431 527 433 703
rect 433 527 485 703
rect 485 527 487 703
rect 115 33 117 209
rect 117 33 169 209
rect 169 33 171 209
rect 273 33 275 209
rect 275 33 327 209
rect 327 33 329 209
<< metal3 >>
rect 105 2082 497 2158
rect 105 1525 181 2082
rect 105 1349 115 1525
rect 171 1349 181 1525
rect 105 209 181 1349
rect 263 1525 339 1530
rect 263 1349 273 1525
rect 329 1349 339 1525
rect 263 1031 339 1349
rect 263 855 273 1031
rect 329 855 339 1031
rect 263 850 339 855
rect 421 1031 497 2082
rect 421 855 431 1031
rect 487 855 497 1031
rect 105 33 115 209
rect 171 33 181 209
rect 105 -524 181 33
rect 263 703 339 708
rect 263 527 273 703
rect 329 527 339 703
rect 263 209 339 527
rect 263 33 273 209
rect 329 33 339 209
rect 263 28 339 33
rect 421 703 497 855
rect 421 527 431 703
rect 487 527 497 703
rect 421 -524 497 527
rect 105 -600 497 -524
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729259347
transform 1 0 99 0 1 943
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729259347
transform 1 0 99 0 1 121
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729259347
transform 1 0 503 0 1 943
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729259347
transform 1 0 503 0 1 615
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729259347
transform 1 0 503 0 1 1437
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729259347
transform 1 0 503 0 1 121
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729259347
transform 1 0 99 0 1 615
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729259347
transform 1 0 99 0 1 1437
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_6HVNUH  sky130_fd_pr__pfet_01v8_6HVNUH_0
timestamp 1729242668
transform 1 0 301 0 1 779
box -223 -364 223 364
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729242668
transform 1 0 301 0 1 121
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729242668
transform 1 0 301 0 1 1437
box -223 -200 223 200
<< labels >>
flabel metal2 303 777 303 777 0 FreeSans 160 0 0 0 d5
port 0 nsew
flabel via1 548 1434 548 1434 0 FreeSans 160 0 0 0 out
port 1 nsew
flabel via2 144 1436 144 1436 0 FreeSans 160 0 0 0 d6
port 2 nsew
flabel via1 219 1108 219 1108 0 FreeSans 160 0 0 0 vip
port 3 nsew
flabel metal1 220 1273 220 1273 0 FreeSans 160 0 0 0 vin
port 4 nsew
flabel viali 303 2173 303 2173 0 FreeSans 160 0 0 0 vdd
port 5 nsew
<< end >>
