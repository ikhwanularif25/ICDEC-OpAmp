magic
tech sky130A
magscale 1 2
timestamp 1729242668
<< nwell >>
rect -325 -483 325 483
<< pmos >>
rect -129 64 -29 264
rect 29 64 129 264
rect -129 -264 -29 -64
rect 29 -264 129 -64
<< pdiff >>
rect -187 252 -129 264
rect -187 76 -175 252
rect -141 76 -129 252
rect -187 64 -129 76
rect -29 252 29 264
rect -29 76 -17 252
rect 17 76 29 252
rect -29 64 29 76
rect 129 252 187 264
rect 129 76 141 252
rect 175 76 187 252
rect 129 64 187 76
rect -187 -76 -129 -64
rect -187 -252 -175 -76
rect -141 -252 -129 -76
rect -187 -264 -129 -252
rect -29 -76 29 -64
rect -29 -252 -17 -76
rect 17 -252 29 -76
rect -29 -264 29 -252
rect 129 -76 187 -64
rect 129 -252 141 -76
rect 175 -252 187 -76
rect 129 -264 187 -252
<< pdiffc >>
rect -175 76 -141 252
rect -17 76 17 252
rect 141 76 175 252
rect -175 -252 -141 -76
rect -17 -252 17 -76
rect 141 -252 175 -76
<< nsubdiff >>
rect -289 413 -193 447
rect 193 413 289 447
rect -289 351 -255 413
rect 255 351 289 413
rect -289 -413 -255 -351
rect 255 -413 289 -351
rect -289 -447 -193 -413
rect 193 -447 289 -413
<< nsubdiffcont >>
rect -193 413 193 447
rect -289 -351 -255 351
rect 255 -351 289 351
rect -193 -447 193 -413
<< poly >>
rect -129 345 -29 361
rect -129 311 -113 345
rect -45 311 -29 345
rect -129 264 -29 311
rect 29 345 129 361
rect 29 311 45 345
rect 113 311 129 345
rect 29 264 129 311
rect -129 17 -29 64
rect -129 -17 -113 17
rect -45 -17 -29 17
rect -129 -64 -29 -17
rect 29 17 129 64
rect 29 -17 45 17
rect 113 -17 129 17
rect 29 -64 129 -17
rect -129 -311 -29 -264
rect -129 -345 -113 -311
rect -45 -345 -29 -311
rect -129 -361 -29 -345
rect 29 -311 129 -264
rect 29 -345 45 -311
rect 113 -345 129 -311
rect 29 -361 129 -345
<< polycont >>
rect -113 311 -45 345
rect 45 311 113 345
rect -113 -17 -45 17
rect 45 -17 113 17
rect -113 -345 -45 -311
rect 45 -345 113 -311
<< locali >>
rect -289 413 -193 447
rect 193 413 289 447
rect -289 351 -255 413
rect 255 351 289 413
rect -129 311 -113 345
rect -45 311 -29 345
rect 29 311 45 345
rect 113 311 129 345
rect -175 252 -141 268
rect -175 60 -141 76
rect -17 252 17 268
rect -17 60 17 76
rect 141 252 175 268
rect 141 60 175 76
rect -129 -17 -113 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 113 -17 129 17
rect -175 -76 -141 -60
rect -175 -268 -141 -252
rect -17 -76 17 -60
rect -17 -268 17 -252
rect 141 -76 175 -60
rect 141 -268 175 -252
rect -129 -345 -113 -311
rect -45 -345 -29 -311
rect 29 -345 45 -311
rect 113 -345 129 -311
rect -289 -413 -255 -351
rect 255 -413 289 -351
rect -289 -447 -193 -413
rect 193 -447 289 -413
<< viali >>
rect -113 311 -45 345
rect 45 311 113 345
rect -175 76 -141 252
rect -17 76 17 252
rect 141 76 175 252
rect -113 -17 -45 17
rect 45 -17 113 17
rect -175 -252 -141 -76
rect -17 -252 17 -76
rect 141 -252 175 -76
rect -113 -345 -45 -311
rect 45 -345 113 -311
<< metal1 >>
rect -125 345 -33 351
rect -125 311 -113 345
rect -45 311 -33 345
rect -125 305 -33 311
rect 33 345 125 351
rect 33 311 45 345
rect 113 311 125 345
rect 33 305 125 311
rect -181 252 -135 264
rect -181 76 -175 252
rect -141 76 -135 252
rect -181 64 -135 76
rect -23 252 23 264
rect -23 76 -17 252
rect 17 76 23 252
rect -23 64 23 76
rect 135 252 181 264
rect 135 76 141 252
rect 175 76 181 252
rect 135 64 181 76
rect -125 17 -33 23
rect -125 -17 -113 17
rect -45 -17 -33 17
rect -125 -23 -33 -17
rect 33 17 125 23
rect 33 -17 45 17
rect 113 -17 125 17
rect 33 -23 125 -17
rect -181 -76 -135 -64
rect -181 -252 -175 -76
rect -141 -252 -135 -76
rect -181 -264 -135 -252
rect -23 -76 23 -64
rect -23 -252 -17 -76
rect 17 -252 23 -76
rect -23 -264 23 -252
rect 135 -76 181 -64
rect 135 -252 141 -76
rect 175 -252 181 -76
rect 135 -264 181 -252
rect -125 -311 -33 -305
rect -125 -345 -113 -311
rect -45 -345 -33 -311
rect -125 -351 -33 -345
rect 33 -311 125 -305
rect 33 -345 45 -311
rect 113 -345 125 -311
rect 33 -351 125 -345
<< properties >>
string FIXED_BBOX -272 -430 272 430
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
