magic
tech sky130A
magscale 1 2
timestamp 1729231875
<< nmos >>
rect -407 55 -247 255
rect -189 55 -29 255
rect 29 55 189 255
rect 247 55 407 255
rect -407 -255 -247 -55
rect -189 -255 -29 -55
rect 29 -255 189 -55
rect 247 -255 407 -55
<< ndiff >>
rect -465 243 -407 255
rect -465 67 -453 243
rect -419 67 -407 243
rect -465 55 -407 67
rect -247 243 -189 255
rect -247 67 -235 243
rect -201 67 -189 243
rect -247 55 -189 67
rect -29 243 29 255
rect -29 67 -17 243
rect 17 67 29 243
rect -29 55 29 67
rect 189 243 247 255
rect 189 67 201 243
rect 235 67 247 243
rect 189 55 247 67
rect 407 243 465 255
rect 407 67 419 243
rect 453 67 465 243
rect 407 55 465 67
rect -465 -67 -407 -55
rect -465 -243 -453 -67
rect -419 -243 -407 -67
rect -465 -255 -407 -243
rect -247 -67 -189 -55
rect -247 -243 -235 -67
rect -201 -243 -189 -67
rect -247 -255 -189 -243
rect -29 -67 29 -55
rect -29 -243 -17 -67
rect 17 -243 29 -67
rect -29 -255 29 -243
rect 189 -67 247 -55
rect 189 -243 201 -67
rect 235 -243 247 -67
rect 189 -255 247 -243
rect 407 -67 465 -55
rect 407 -243 419 -67
rect 453 -243 465 -67
rect 407 -255 465 -243
<< ndiffc >>
rect -453 67 -419 243
rect -235 67 -201 243
rect -17 67 17 243
rect 201 67 235 243
rect 419 67 453 243
rect -453 -243 -419 -67
rect -235 -243 -201 -67
rect -17 -243 17 -67
rect 201 -243 235 -67
rect 419 -243 453 -67
<< poly >>
rect -407 327 -247 343
rect -407 293 -391 327
rect -263 293 -247 327
rect -407 255 -247 293
rect -189 327 -29 343
rect -189 293 -173 327
rect -45 293 -29 327
rect -189 255 -29 293
rect 29 327 189 343
rect 29 293 45 327
rect 173 293 189 327
rect 29 255 189 293
rect 247 327 407 343
rect 247 293 263 327
rect 391 293 407 327
rect 247 255 407 293
rect -407 17 -247 55
rect -407 -17 -391 17
rect -263 -17 -247 17
rect -407 -55 -247 -17
rect -189 17 -29 55
rect -189 -17 -173 17
rect -45 -17 -29 17
rect -189 -55 -29 -17
rect 29 17 189 55
rect 29 -17 45 17
rect 173 -17 189 17
rect 29 -55 189 -17
rect 247 17 407 55
rect 247 -17 263 17
rect 391 -17 407 17
rect 247 -55 407 -17
rect -407 -293 -247 -255
rect -407 -327 -391 -293
rect -263 -327 -247 -293
rect -407 -343 -247 -327
rect -189 -293 -29 -255
rect -189 -327 -173 -293
rect -45 -327 -29 -293
rect -189 -343 -29 -327
rect 29 -293 189 -255
rect 29 -327 45 -293
rect 173 -327 189 -293
rect 29 -343 189 -327
rect 247 -293 407 -255
rect 247 -327 263 -293
rect 391 -327 407 -293
rect 247 -343 407 -327
<< polycont >>
rect -391 293 -263 327
rect -173 293 -45 327
rect 45 293 173 327
rect 263 293 391 327
rect -391 -17 -263 17
rect -173 -17 -45 17
rect 45 -17 173 17
rect 263 -17 391 17
rect -391 -327 -263 -293
rect -173 -327 -45 -293
rect 45 -327 173 -293
rect 263 -327 391 -293
<< locali >>
rect -407 293 -391 327
rect -263 293 -247 327
rect -189 293 -173 327
rect -45 293 -29 327
rect 29 293 45 327
rect 173 293 189 327
rect 247 293 263 327
rect 391 293 407 327
rect -453 243 -419 259
rect -453 51 -419 67
rect -235 243 -201 259
rect -235 51 -201 67
rect -17 243 17 259
rect -17 51 17 67
rect 201 243 235 259
rect 201 51 235 67
rect 419 243 453 259
rect 419 51 453 67
rect -407 -17 -391 17
rect -263 -17 -247 17
rect -189 -17 -173 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 173 -17 189 17
rect 247 -17 263 17
rect 391 -17 407 17
rect -453 -67 -419 -51
rect -453 -259 -419 -243
rect -235 -67 -201 -51
rect -235 -259 -201 -243
rect -17 -67 17 -51
rect -17 -259 17 -243
rect 201 -67 235 -51
rect 201 -259 235 -243
rect 419 -67 453 -51
rect 419 -259 453 -243
rect -407 -327 -391 -293
rect -263 -327 -247 -293
rect -189 -327 -173 -293
rect -45 -327 -29 -293
rect 29 -327 45 -293
rect 173 -327 189 -293
rect 247 -327 263 -293
rect 391 -327 407 -293
<< viali >>
rect -391 293 -263 327
rect -173 293 -45 327
rect 45 293 173 327
rect 263 293 391 327
rect -453 67 -419 243
rect -235 67 -201 243
rect -17 67 17 243
rect 201 67 235 243
rect 419 67 453 243
rect -391 -17 -263 17
rect -173 -17 -45 17
rect 45 -17 173 17
rect 263 -17 391 17
rect -453 -243 -419 -67
rect -235 -243 -201 -67
rect -17 -243 17 -67
rect 201 -243 235 -67
rect 419 -243 453 -67
rect -391 -327 -263 -293
rect -173 -327 -45 -293
rect 45 -327 173 -293
rect 263 -327 391 -293
<< metal1 >>
rect -403 327 -251 333
rect -403 293 -391 327
rect -263 293 -251 327
rect -403 287 -251 293
rect -185 327 -33 333
rect -185 293 -173 327
rect -45 293 -33 327
rect -185 287 -33 293
rect 33 327 185 333
rect 33 293 45 327
rect 173 293 185 327
rect 33 287 185 293
rect 251 327 403 333
rect 251 293 263 327
rect 391 293 403 327
rect 251 287 403 293
rect -459 243 -413 255
rect -459 67 -453 243
rect -419 67 -413 243
rect -459 55 -413 67
rect -241 243 -195 255
rect -241 67 -235 243
rect -201 67 -195 243
rect -241 55 -195 67
rect -23 243 23 255
rect -23 67 -17 243
rect 17 67 23 243
rect -23 55 23 67
rect 195 243 241 255
rect 195 67 201 243
rect 235 67 241 243
rect 195 55 241 67
rect 413 243 459 255
rect 413 67 419 243
rect 453 67 459 243
rect 413 55 459 67
rect -403 17 -251 23
rect -403 -17 -391 17
rect -263 -17 -251 17
rect -403 -23 -251 -17
rect -185 17 -33 23
rect -185 -17 -173 17
rect -45 -17 -33 17
rect -185 -23 -33 -17
rect 33 17 185 23
rect 33 -17 45 17
rect 173 -17 185 17
rect 33 -23 185 -17
rect 251 17 403 23
rect 251 -17 263 17
rect 391 -17 403 17
rect 251 -23 403 -17
rect -459 -67 -413 -55
rect -459 -243 -453 -67
rect -419 -243 -413 -67
rect -459 -255 -413 -243
rect -241 -67 -195 -55
rect -241 -243 -235 -67
rect -201 -243 -195 -67
rect -241 -255 -195 -243
rect -23 -67 23 -55
rect -23 -243 -17 -67
rect 17 -243 23 -67
rect -23 -255 23 -243
rect 195 -67 241 -55
rect 195 -243 201 -67
rect 235 -243 241 -67
rect 195 -255 241 -243
rect 413 -67 459 -55
rect 413 -243 419 -67
rect 453 -243 459 -67
rect 413 -255 459 -243
rect -403 -293 -251 -287
rect -403 -327 -391 -293
rect -263 -327 -251 -293
rect -403 -333 -251 -327
rect -185 -293 -33 -287
rect -185 -327 -173 -293
rect -45 -327 -33 -293
rect -185 -333 -33 -327
rect 33 -293 185 -287
rect 33 -327 45 -293
rect 173 -327 185 -293
rect 33 -333 185 -327
rect 251 -293 403 -287
rect 251 -327 263 -293
rect 391 -327 403 -293
rect 251 -333 403 -327
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
