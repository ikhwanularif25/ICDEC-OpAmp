magic
tech sky130A
magscale 1 2
timestamp 1729158022
<< nmos >>
rect -229 -231 -29 169
rect 29 -231 229 169
<< ndiff >>
rect -287 157 -229 169
rect -287 -219 -275 157
rect -241 -219 -229 157
rect -287 -231 -229 -219
rect -29 157 29 169
rect -29 -219 -17 157
rect 17 -219 29 157
rect -29 -231 29 -219
rect 229 157 287 169
rect 229 -219 241 157
rect 275 -219 287 157
rect 229 -231 287 -219
<< ndiffc >>
rect -275 -219 -241 157
rect -17 -219 17 157
rect 241 -219 275 157
<< poly >>
rect -229 241 -29 257
rect -229 207 -213 241
rect -45 207 -29 241
rect -229 169 -29 207
rect 29 241 229 257
rect 29 207 45 241
rect 213 207 229 241
rect 29 169 229 207
rect -229 -257 -29 -231
rect 29 -257 229 -231
<< polycont >>
rect -213 207 -45 241
rect 45 207 213 241
<< locali >>
rect -229 207 -213 241
rect -45 207 -29 241
rect 29 207 45 241
rect 213 207 229 241
rect -275 157 -241 173
rect -275 -235 -241 -219
rect -17 157 17 173
rect -17 -235 17 -219
rect 241 157 275 173
rect 241 -235 275 -219
<< viali >>
rect -213 207 -45 241
rect 45 207 213 241
rect -275 -219 -241 157
rect -17 -219 17 157
rect 241 -219 275 157
<< metal1 >>
rect -225 241 -33 247
rect -225 207 -213 241
rect -45 207 -33 241
rect -225 201 -33 207
rect 33 241 225 247
rect 33 207 45 241
rect 213 207 225 241
rect 33 201 225 207
rect -281 157 -235 169
rect -281 -219 -275 157
rect -241 -219 -235 157
rect -281 -231 -235 -219
rect -23 157 23 169
rect -23 -219 -17 157
rect 17 -219 23 157
rect -23 -231 23 -219
rect 235 157 281 169
rect 235 -219 241 157
rect 275 -219 281 157
rect 235 -231 281 -219
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
