magic
tech sky130A
magscale 1 2
timestamp 1729220960
<< error_p >>
rect -29 381 29 387
rect -29 347 -17 381
rect -29 341 29 347
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect -29 -387 29 -381
<< nmos >>
rect -15 109 15 309
rect -15 -309 15 -109
<< ndiff >>
rect -73 297 -15 309
rect -73 121 -61 297
rect -27 121 -15 297
rect -73 109 -15 121
rect 15 297 73 309
rect 15 121 27 297
rect 61 121 73 297
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -297 -61 -121
rect -27 -297 -15 -121
rect -73 -309 -15 -297
rect 15 -121 73 -109
rect 15 -297 27 -121
rect 61 -297 73 -121
rect 15 -309 73 -297
<< ndiffc >>
rect -61 121 -27 297
rect 27 121 61 297
rect -61 -297 -27 -121
rect 27 -297 61 -121
<< poly >>
rect -33 381 33 397
rect -33 347 -17 381
rect 17 347 33 381
rect -33 331 33 347
rect -15 309 15 331
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -331 15 -309
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
<< polycont >>
rect -17 347 17 381
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -381 17 -347
<< locali >>
rect -33 347 -17 381
rect 17 347 33 381
rect -61 297 -27 313
rect -61 105 -27 121
rect 27 297 61 313
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -313 -27 -297
rect 27 -121 61 -105
rect 27 -313 61 -297
rect -33 -381 -17 -347
rect 17 -381 33 -347
<< viali >>
rect -17 347 17 381
rect -61 121 -27 297
rect 27 121 61 297
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -297 -27 -121
rect 27 -297 61 -121
rect -17 -381 17 -347
<< metal1 >>
rect -29 381 29 387
rect -29 347 -17 381
rect 17 347 29 381
rect -29 341 29 347
rect -67 297 -21 309
rect -67 121 -61 297
rect -27 121 -21 297
rect -67 109 -21 121
rect 21 297 67 309
rect 21 121 27 297
rect 61 121 67 297
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -297 -61 -121
rect -27 -297 -21 -121
rect -67 -309 -21 -297
rect 21 -121 67 -109
rect 21 -297 27 -121
rect 61 -297 67 -121
rect 21 -309 67 -297
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
